module main

import term.ui as tui

const color_black = tui.Color{
	r: 0
	g: 0
	b: 0
}
const color_green = tui.Color{
	r: 0
	g: 228
	b: 54
}
const color_blue = tui.Color{
	r: 41
	g: 173
	b: 255
}
const color_yellow = tui.Color{
	r: 255
	g: 236
	b: 39
}
const color_red = tui.Color{
	r: 255
	g: 0
	b: 77
}
